// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_proj_example
 *
 * This is an example of a (trivially simple) user project,
 * showing how the user project can connect to the logic
 * analyzer, the wishbone bus, and the I/O pads.
 *
 * This project generates an integer count, which is output
 * on the user area GPIO pads (digital output only).  The
 * wishbone connection allows the project to be controlled
 * (start and stop) from the management SoC program.
 *
 * See the testbenches in directory "mprj_counter" for the
 * example programs that drive this user project.  The three
 * testbenches are "io_ports", "la_test1", and "la_test2".
 *
 *-------------------------------------------------------------
 */

module user_proj_example #(
    parameter BITS = 32
)(
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // IRQ
    output [2:0] irq
);
    wire clk;
    wire rst;

    wire [`MPRJ_IO_PADS-1:0] io_in;
    wire [`MPRJ_IO_PADS-1:0] io_out;
    wire [`MPRJ_IO_PADS-1:0] io_oeb;

    wire [31:0] rdata; 
    wire [31:0] wdata;
    wire [BITS-1:0] count;

    wire valid;
    wire [3:0] wstrb;
    wire [31:0] la_write;

    // WB MI A
    assign valid = wbs_cyc_i && wbs_stb_i; 
    assign wstrb = wbs_sel_i & {4{wbs_we_i}};
    assign wbs_dat_o = rdata;
    assign wdata = wbs_dat_i;

    // IO
    assign io_out = count;
    assign io_oeb = {(`MPRJ_IO_PADS-1){rst}};

    // IRQ
    assign irq = 3'b000;	// Unused

    // LA
    assign la_data_out = {{(127-BITS){1'b0}}, count};
    // Assuming LA probes [63:32] are for controlling the count register  
    assign la_write = ~la_oenb[63:32] & ~{BITS{valid}};
    // Assuming LA probes [65:64] are for controlling the count clk & reset  
    assign clk = (~la_oenb[64]) ? la_data_in[64]: wb_clk_i;
    assign rst = (~la_oenb[65]) ? la_data_in[65]: wb_rst_i;

pro_row_idct_parallel dut(

i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
s,se,

ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,

ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,

ou80s,ou81s,ou82s,ou83s,
ou80,ou81,ou82,ou83,

ou160s,ou161s,
ou160,ou161,

ou320s,
ou320

);


endmodule

//proposed 32-point configurable IntegerDCT for row process in parallel architecture

//`include "block_complete_row_parallel.v"
////`include "cell_sign.v"
//`include "adder24.v"

module pro_row_idct_parallel(

i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,
i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
s,se,

ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,

ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,

ou80s,ou81s,ou82s,ou83s,
ou80,ou81,ou82,ou83,

ou160s,ou161s,
ou160,ou161,

ou320s,
ou320

);

output ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou80s,ou81s,ou82s,ou83s,
ou160s,ou161s,
ou320s;

output [23:0] ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,
ou80,ou81,ou82,ou83,
ou160,ou161,
ou320;

input i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s;
input [7:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31;

input [4:0] s;
input [2:0] se;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

wire [23:0] o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,o20,o21,o22,o23,o24,o25,o26,o27,o28,o29,o30,o31;
wire o0s,o1s,o2s,o3s,o4s,o5s,o6s,o7s,o8s,o9s,o10s,o11s,o12s,o13s,o14s,o15s,o16s,o17s,o18s,o19s,o20s,o21s,o22s,o23s,o24s,o25s,o26s,o27s,o28s,o29s,o30s,o31s;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp0(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o0

);

cell_sign cc0(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o0s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp1(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o1

);

cell_sign cc1(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o1s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp2(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o2

);

cell_sign cc2(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o2s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp3(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o3

);

cell_sign cc3(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o3s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp4(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o4

);

cell_sign cc4(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o4s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp5(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o5

);

cell_sign cc5(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o5s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp6(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o6

);

cell_sign cc6(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o6s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp7(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o7

);

cell_sign cc7(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o7s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp8(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o8

);

cell_sign cc8(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o8s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp9(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o9

);

cell_sign cc9(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o9s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp10(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o10

);

cell_sign cc10(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o10s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp11(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o11

);

cell_sign cc11(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o11s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp12(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o12

);

cell_sign cc12(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o12s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp13(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o13

);

cell_sign cc13(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o13s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp14(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o14

);

cell_sign cc14(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o14s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp15(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o15

);

cell_sign cc15(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o15s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp16(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o16

);

cell_sign cc16(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o16s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp17(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o17

);

cell_sign cc17(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o17s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp18(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o18

);

cell_sign cc18(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o18s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp19(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o19

);

cell_sign cc19(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o19s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp20(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o20

);

cell_sign cc20(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o20s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp21(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o21

);

cell_sign cc21(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o21s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp22(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o22

);

cell_sign cc22(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o22s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp23(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o23

);

cell_sign cc23(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o23s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp24(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o24

);

cell_sign cc24(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o24s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp25(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o25

);

cell_sign cc25(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o25s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp26(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o26

);

cell_sign cc26(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o26s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp27(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o27

);

cell_sign cc27(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o27s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp28(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o28

);

cell_sign cc28(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o28s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp29(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o29

);

cell_sign cc29(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o29s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp30(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o30

);

cell_sign cc30(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o30s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

block_complete_row_parallel pp31(

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},{16'd0,i16},{16'd0,i17},{16'd0,i18},{16'd0,i19},{16'd0,i20},{16'd0,i21},{16'd0,i22},{16'd0,i23},{16'd0,i24},{16'd0,i25},{16'd0,i26},{16'd0,i27},{16'd0,i28},{16'd0,i29},{16'd0,i30},{16'd0,i31},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},{16'd0,i8},{16'd0,i9},{16'd0,i10},{16'd0,i11},{16'd0,i12},{16'd0,i13},{16'd0,i14},{16'd0,i15},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},{16'd0,i4},{16'd0,i5},{16'd0,i6},{16'd0,i7},
{16'd0,i0},{16'd0,i1},{16'd0,i2},{16'd0,i3},
{16'd0,i0},{16'd0,i1},

s,se,o31

);

cell_sign cc31(i0s,i1s,i2s,i3s,i4s,i5s,i6s,i7s,i8s,i9s,i10s,i11s,i12s,i13s,i14s,i15s,i16s,i17s,i18s,i19s,i20s,i21s,i22s,i23s,i24s,i25s,i26s,i27s,i28s,i29s,i30s,i31s,s,se,o31s);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

wire ou20s,ou21s,ou22s,ou23s,ou24s,ou25s,ou26s,ou27s,ou28s,ou29s,ou210s,ou211s,ou212s,ou213s,ou214s,ou215s,
ou40s,ou41s,ou42s,ou43s,ou44s,ou45s,ou46s,ou47s,
ou80s,ou81s,ou82s,ou83s,
ou160s,ou161s,
ou320s;

wire [23:0] ou20,ou21,ou22,ou23,ou24,ou25,ou26,ou27,ou28,ou29,ou210,ou211,ou212,ou213,ou214,ou215,
ou40,ou41,ou42,ou43,ou44,ou45,ou46,ou47,
ou80,ou81,ou82,ou83,
ou160,ou161,
ou320;

//first level of tree of adders

adder24 ad10(o0s,o0,o1s,o1,ou20s,ou20);
adder24 ad11(o2s,o2,o3s,o3,ou21s,ou21);
adder24 ad12(o4s,o4,o5s,o5,ou22s,ou22);
adder24 ad13(o6s,o6,o7s,o7,ou23s,ou23);
adder24 ad14(o8s,o8,o9s,o9,ou24s,ou24);
adder24 ad15(o10s,o10,o11s,o11,ou25s,ou25);
adder24 ad16(o12s,o12,o13s,o13,ou26s,ou26);
adder24 ad17(o14s,o14,o15s,o15,ou27s,ou27);
adder24 ad18(o16s,o16,o17s,o17,ou28s,ou28);
adder24 ad19(o18s,o18,o19s,o19,ou29s,ou29);
adder24 ad110(o20s,o20,o21s,o21,ou210s,ou210);
adder24 ad111(o22s,o22,o23s,o23,ou211s,ou211);
adder24 ad112(o24s,o24,o25s,o25,ou212s,ou212);
adder24 ad113(o26s,o26,o27s,o27,ou213s,ou213);
adder24 ad114(o28s,o28,o29s,o29,ou214s,ou214);
adder24 ad115(o30s,o30,o31s,o31,ou215s,ou215);

//second level of tree of adders

adder24 ad20(ou20s,ou20,ou21s,ou21,ou40s,ou40);
adder24 ad21(ou22s,ou22,ou23s,ou23,ou41s,ou41);
adder24 ad22(ou24s,ou24,ou25s,ou25,ou42s,ou42);
adder24 ad23(ou26s,ou26,ou27s,ou27,ou43s,ou43);
adder24 ad24(ou28s,ou28,ou29s,ou29,ou44s,ou44);
adder24 ad25(ou210s,ou210,ou211s,ou211,ou45s,ou45);
adder24 ad26(ou212s,ou212,ou213s,ou213,ou46s,ou46);
adder24 ad27(ou214s,ou214,ou215s,ou215,ou47s,ou47);

//third level of tree of adders

adder24 ad30(ou40s,ou40,ou41s,ou41,ou80s,ou80);
adder24 ad31(ou42s,ou42,ou43s,ou43,ou81s,ou81);
adder24 ad32(ou44s,ou44,ou45s,ou45,ou82s,ou82);
adder24 ad33(ou46s,ou46,ou47s,ou47,ou83s,ou83);

//fourth level of tree of adders

adder24 ad40(ou80s,ou80,ou81s,ou81,ou160s,ou160);
adder24 ad41(ou82s,ou82,ou83s,ou83,ou161s,ou161);

//fifth level of tree of adders

adder24 ad50(ou160s,ou160,ou161s,ou161,ou320s,ou320);

endmodule


//24 bit fixed point adder

//`include "recurse24.v"
//`include "kgp.v"
//`include "kgp_carry.v"
//`include "recursive_stage1.v"

module adder24(as,a,bs,in_b,rrs,rr);

input as,bs;
input [23:0] a,in_b;
output rrs;
output [23:0] rr;

reg rrs;
reg [23:0] rr;
wire z;
assign z=as^bs;
wire cout,cout1;

wire [23:0] r1,b1,b2;
assign b1=(~in_b);

recurse24 c0(b2,cout1,b1,24'b000000000000000000000001);

reg [23:0] b;

always@(z or in_b or b2)
	begin
		if(z==0)
			b=in_b;
		else if (z==1)
			b=b2;
	end
	
recurse24 c1(r1,cout,a,b);

wire cout2;
wire [23:0] r11,r22;
assign r11=(~r1);
recurse24 c2(r22,cout2,r11,24'b000000000000000000000001);

reg carry;
always@(r1 or cout or z or as or bs or r22)
 begin
	if(z==0)	
		begin
			rrs=as;
			rr=r1;
			carry=cout;
		end
	else if (z==1 && cout==1)
		begin	
			rrs=as;
			rr=r1;
			carry=1'b0;
		end
	else if (z==1 && cout==0)
		begin
			rrs=(~as);
			rr=r22;
			carry=1'b0;
		end
 end

endmodule


/*`include "mux32to1_1.v"
`include "mux16to1_1.v"
`include "mux8to1_1.v"
`include "mux4to1_1.v"
`include "mux2to1_1.v"
`include "mux5to1_1.v"*/

//cell used for sign in Integer DCT 

module cell_sign(i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,s,se,out);

input i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31;
input [4:0] s;
input [2:0] se;
output out;

wire out1,out2,out3,out4,out5;

wire si0,si1,si2,si3,si4,si5,si6,si7,si8,si9,si10,si11,si12,si13,si14,si15,si16,si17,si18,si19,si20,si21,si22,si23,si24,si25,si26,si27,si28,si29,si30,si31;

assign si0=i0^1'b0;
assign si1=i1^1'b0;
assign si2=i2^1'b0;
assign si3=i3^1'b0;
assign si4=i4^1'b0;
assign si5=i5^1'b0;
assign si6=i6^1'b0;
assign si7=i7^1'b0;
assign si8=i8^1'b0;
assign si9=i9^1'b0;
assign si10=i10^1'b0;
assign si11=i11^1'b0;
assign si12=i12^1'b0;
assign si13=i13^1'b0;
assign si14=i14^1'b0;
assign si15=i15^1'b0;
assign si16=i16^1'b0;
assign si17=i17^1'b0;
assign si18=i18^1'b0;
assign si19=i19^1'b0;
assign si20=i20^1'b0;
assign si21=i21^1'b0;
assign si22=i22^1'b0;
assign si23=i23^1'b0;
assign si24=i24^1'b0;
assign si25=i25^1'b0;
assign si26=i26^1'b0;
assign si27=i27^1'b0;
assign si28=i28^1'b0;
assign si29=i29^1'b0;
assign si30=i30^1'b0;
assign si31=i31^1'b0;

mux32to1_1 mu1(out1,si0,si1,si2,si3,si4,si5,si6,si7,si8,si9,si10,si11,si12,si13,si14,si15,si16,si17,si18,si19,si20,si21,si22,si23,si24,si25,si26,si27,si28,si29,si30,si31,s[4],s[3],s[2],s[1],s[0]);
mux16to1_1 mu2(out2,si0,si1,si2,si3,si4,si5,si6,si7,si8,si9,si10,si11,si12,si13,si14,si15,s[3:0]);
mux8to1_1 mmu3(out3,si0,si1,si2,si3,si4,si5,si6,si7,s[2:0]);
mux4to1_1 mmu4(out4,si0,si1,si2,si3,s[1:0]);
mux2to1_1 mmu5(out5,si0,si1,s[0]);
mux5to1_1 mmu6(out,out1,out2,out3,out4,out5,se);

endmodule



//The complete block used for row process in parallel architecture

//`include "cell_row_parallel.v"
//`include "block_row_parallel.v"

module block_complete_row_parallel(

i00,i01,i02,i03,i04,i05,i06,i07,i08,i09,i010,i011,i012,i013,i014,i015,i016,i017,i018,i019,i020,i021,i022,i023,i024,i025,i026,i027,i028,i029,i030,i031,
n00,n01,n02,n03,n04,n05,n06,n07,n08,n09,n010,n011,n012,n013,n014,n015,
m00,m01,m02,m03,m04,m05,m06,m07,
o00,o01,o02,o03,
p00,p01,

i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,i130,i131,
n10,n11,n12,n13,n14,n15,n16,n17,n18,n19,n110,n111,n112,n113,n114,n115,
m10,m11,m12,m13,m14,m15,m16,m17,
o10,o11,o12,o13,
p10,p11,

i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i210,i211,i212,i213,i214,i215,i216,i217,i218,i219,i220,i221,i222,i223,i224,i225,i226,i227,i228,i229,i230,i231,
n20,n21,n22,n23,n24,n25,n26,n27,n28,n29,n210,n211,n212,n213,n214,n215,
m20,m21,m22,m23,m24,m25,m26,m27,
o20,o21,o22,o23,
p20,p21,

i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,i310,i311,i312,i313,i314,i315,i316,i317,i318,i319,i320,i321,i322,i323,i324,i325,i326,i327,i328,i329,i330,i331,
n30,n31,n32,n33,n34,n35,n36,n37,n38,n39,n310,n311,n312,n313,n314,n315,
m30,m31,m32,m33,m34,m35,m36,m37,
o30,o31,o32,o33,
p30,p31,

i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,i410,i411,i412,i413,i414,i415,i416,i417,i418,i419,i420,i421,i422,i423,i424,i425,i426,i427,i428,i429,i430,i431,
n40,n41,n42,n43,n44,n45,n46,n47,n48,n49,n410,n411,n412,n413,n414,n415,
m40,m41,m42,m43,m44,m45,m46,m47,
o40,o41,o42,o43,
p40,p41,

s,se,out

);

output [23:0] out;

input [4:0] s;
input [2:0] se;

input [23:0] i00,i01,i02,i03,i04,i05,i06,i07,i08,i09,i010,i011,i012,i013,i014,i015,i016,i017,i018,i019,i020,i021,i022,i023,i024,i025,i026,i027,i028,i029,i030,i031,
n00,n01,n02,n03,n04,n05,n06,n07,n08,n09,n010,n011,n012,n013,n014,n015,
m00,m01,m02,m03,m04,m05,m06,m07,
o00,o01,o02,o03,
p00,p01,

i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,i130,i131,
n10,n11,n12,n13,n14,n15,n16,n17,n18,n19,n110,n111,n112,n113,n114,n115,
m10,m11,m12,m13,m14,m15,m16,m17,
o10,o11,o12,o13,
p10,p11,

i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i210,i211,i212,i213,i214,i215,i216,i217,i218,i219,i220,i221,i222,i223,i224,i225,i226,i227,i228,i229,i230,i231,
n20,n21,n22,n23,n24,n25,n26,n27,n28,n29,n210,n211,n212,n213,n214,n215,
m20,m21,m22,m23,m24,m25,m26,m27,
o20,o21,o22,o23,
p20,p21,

i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,i310,i311,i312,i313,i314,i315,i316,i317,i318,i319,i320,i321,i322,i323,i324,i325,i326,i327,i328,i329,i330,i331,
n30,n31,n32,n33,n34,n35,n36,n37,n38,n39,n310,n311,n312,n313,n314,n315,
m30,m31,m32,m33,m34,m35,m36,m37,
o30,o31,o32,o33,
p30,p31,

i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,i410,i411,i412,i413,i414,i415,i416,i417,i418,i419,i420,i421,i422,i423,i424,i425,i426,i427,i428,i429,i430,i431,
n40,n41,n42,n43,n44,n45,n46,n47,n48,n49,n410,n411,n412,n413,n414,n415,
m40,m41,m42,m43,m44,m45,m46,m47,
o40,o41,o42,o43,
p40,p41;

wire [23:0] b0,b1,b2,b3,b4;

cell_row_parallel c0(i00,i01,i02,i03,i04,i05,i06,i07,i08,i09,i010,i011,i012,i013,i014,i015,i016,i017,i018,i019,i020,i021,i022,i023,i024,i025,i026,i027,i028,i029,i030,i031,
n00,n01,n02,n03,n04,n05,n06,n07,n08,n09,n010,n011,n012,n013,n014,n015,
m00,m01,m02,m03,m04,m05,m06,m07,
o00,o01,o02,o03,
p00,p01,
s,se,b0

);

cell_row_parallel c1(i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,i130,i131,
n10,n11,n12,n13,n14,n15,n16,n17,n18,n19,n110,n111,n112,n113,n114,n115,
m10,m11,m12,m13,m14,m15,m16,m17,
o10,o11,o12,o13,
p10,p11,
s,se,b1

);

cell_row_parallel c2(i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i210,i211,i212,i213,i214,i215,i216,i217,i218,i219,i220,i221,i222,i223,i224,i225,i226,i227,i228,i229,i230,i231,
n20,n21,n22,n23,n24,n25,n26,n27,n28,n29,n210,n211,n212,n213,n214,n215,
m20,m21,m22,m23,m24,m25,m26,m27,
o20,o21,o22,o23,
p20,p21,
s,se,b2

);

cell_row_parallel c3(i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,i310,i311,i312,i313,i314,i315,i316,i317,i318,i319,i320,i321,i322,i323,i324,i325,i326,i327,i328,i329,i330,i331,
n30,n31,n32,n33,n34,n35,n36,n37,n38,n39,n310,n311,n312,n313,n314,n315,
m30,m31,m32,m33,m34,m35,m36,m37,
o30,o31,o32,o33,
p30,p31,
s,se,b3

);

cell_row_parallel c4(i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,i410,i411,i412,i413,i414,i415,i416,i417,i418,i419,i420,i421,i422,i423,i424,i425,i426,i427,i428,i429,i430,i431,
n40,n41,n42,n43,n44,n45,n46,n47,n48,n49,n410,n411,n412,n413,n414,n415,
m40,m41,m42,m43,m44,m45,m46,m47,
o40,o41,o42,o43,
p40,p41,
s,se,b4

);

block_row_parallel block(b0,b1,b2,b3,b4,out);

endmodule



/*`include "mux32to1_24.v"
`include "mux16to1_24.v"
`include "mux8to1_24.v"
`include "mux4to1_24.v"
`include "mux2to1_24.v"
`include "mux5to1_24.v"*/

//cell used for row process in parallel architecture of Integer DCT

module cell_row_parallel(i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
n0,n1,n2,n3,n4,n5,n6,n7,n8,n9,n10,n11,n12,n13,n14,n15,
m0,m1,m2,m3,m4,m5,m6,m7,
o0,o1,o2,o3,
p0,p1,
s,se,out

);

input [23:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,
n0,n1,n2,n3,n4,n5,n6,n7,n8,n9,n10,n11,n12,n13,n14,n15,
m0,m1,m2,m3,m4,m5,m6,m7,
o0,o1,o2,o3,
p0,p1;

input [4:0] s;
input [2:0] se;
output [23:0] out;

wire [23:0] out1,out2,out3,out4,out5;

mux32to1_24 mu1(out1,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,s[4],s[3],s[2],s[1],s[0]);
mux16to1_24 mu2(out2,n0,n1,n2,n3,n4,n5,n6,n7,n8,n9,n10,n11,n12,n13,n14,n15,s[3:0]);
mux8to1_24 mmu3(out3,m0,m1,m2,m3,m4,m5,m6,m7,s[2:0]);
mux4to1_24 mmu4(out4,o0,o1,o2,o3,s[1:0]);
mux2to1_24 mmu5(out5,p0,p1,s[0]);
mux5to1_24 mmu6(out,out1,out2,out3,out4,out5,se);

endmodule





/*`include "halfadd.v"
`include "fulladd.v"
`include "kgp.v"
`include "kgp_carry.v"
`include "recursive_stage1.v"*/
//`include "recurse24.v"

//block used for row process in parallel architecture

module block_row_parallel(i0,i1,i2,i3,i4,out);

input [23:0] i0,i1,i2,i3,i4;
output [23:0] out;

wire [23:0] sum1h,sum11h,sum2h;
wire carry1h,carry11h,carry2h,carry;

recurse24 rr1(sum1h,carry1h,i0,i1);
recurse24 rr2(sum11h,carry11h,i2,i3);
recurse24 rr3(sum2h,carry2h,sum1h,sum11h); 
recurse24 rr4(out,carry,sum2h,i4); 

endmodule




module kgp(a,b,y);

input a,b;
output [1:0] y;
//reg [1:0] y;

//always@(a or b)
//begin
//case({a,b})
//2'b00:y=2'b00;  //kill
//2'b11:y=2'b11;	  //generate
//2'b01:y=2'b01;	//propagate
//2'b10:y=2'b01;  //propagate
//endcase   //y[1]=ab  y[0]=a+b  
//end

assign y[0]=a | b;
assign y[1]=a & b;

endmodule




module kgp_carry(a,b,carry);

input [1:0] a,b;
output carry;
reg carry;

always@(a or b)
begin
case(a)
2'b00:carry=1'b0;  
2'b11:carry=1'b1;
2'b01:carry=b[0];
2'b10:carry=b[0];
default:carry=1'bx;
endcase
end

/*wire carry;

wire f,g;
assign g=a[0] & a[1];
assign f=a[0] ^ a[1];

assign carry=g|(b[0] & f);*/

endmodule




module recursive_stage1(a,b,y);

input [1:0] a,b;
output [1:0] y;

wire [1:0] y;
wire b0;
not n1(b0,b[1]);
wire f,g0,g1;
and a1(f,b[0],b[1]);
and a2(g0,b0,b[0],a[0]);
and a3(g1,b0,b[0],a[1]);

or o1(y[0],f,g0);
or o2(y[1],f,g1);

//reg [1:0] y;
//always@(a or b)
//begin
//case(b)
//2'b00:y=2'b00;  
//2'b11:y=2'b11;
//2'b01:y=a;
//default:y=2'bx;
//endcase
//end

//always@(a or b)
//begin
//if(b==2'b00)
//	y=2'b00;  
//else if (b==2'b11)
//	y=2'b11;
//else if (b==2'b01)
//	y=a;
//end

//wire x;
//assign x=a[0] ^ b[0];
//always@(a or b or x)
//begin
//case(x)
//1'b0:y[0]=b[0];  
//1'b1:y[0]=a[0]; 
//endcase
//end
//
//always@(a or b or x)
//begin
//case(x)
//1'b0:y[1]=b[1];  
//1'b1:y[1]=a[1];
//endcase
//end


//always@(a or b)
//begin
//if (b==2'b00)
//	y=2'b00; 
//else if (b==2'b11)	
//	y=2'b11;
//else if (b==2'b01 && a==2'b00)
//	y=2'b00;
//else if (b==2'b01 && a==2'b11)
//	y=2'b11;
//else if (b==2'b01 && a==2'b01)
//	y=2'b01;
//end

endmodule


//24 bit recursive doubling technique

module recurse24(sum,carry,a,b); 

output [23:0] sum;
output  carry;
input [23:0] a,b;

wire [49:0] x;

assign x[1:0]=2'b00;  // kgp generation

kgp a00(a[0],b[0],x[3:2]);
kgp a01(a[1],b[1],x[5:4]);
kgp a02(a[2],b[2],x[7:6]);
kgp a03(a[3],b[3],x[9:8]);
kgp a04(a[4],b[4],x[11:10]);
kgp a05(a[5],b[5],x[13:12]);
kgp a06(a[6],b[6],x[15:14]);
kgp a07(a[7],b[7],x[17:16]);
kgp a08(a[8],b[8],x[19:18]);
kgp a09(a[9],b[9],x[21:20]);
kgp a10(a[10],b[10],x[23:22]);
kgp a11(a[11],b[11],x[25:24]);
kgp a12(a[12],b[12],x[27:26]);
kgp a13(a[13],b[13],x[29:28]);
kgp a14(a[14],b[14],x[31:30]);
kgp a15(a[15],b[15],x[33:32]);
kgp a16(a[16],b[16],x[35:34]);
kgp a17(a[17],b[17],x[37:36]);
kgp a18(a[18],b[18],x[39:38]);
kgp a19(a[19],b[19],x[41:40]);
kgp a20(a[20],b[20],x[43:42]);
kgp a21(a[21],b[21],x[45:44]);
kgp a22(a[22],b[22],x[47:46]);
kgp a23(a[23],b[23],x[49:48]);

wire [49:0] x1;  //recursive doubling stage 1
assign x1[1:0]=x[1:0];

recursive_stage1 s00(x[1:0],x[3:2],x1[3:2]);
recursive_stage1 s01(x[3:2],x[5:4],x1[5:4]);
recursive_stage1 s02(x[5:4],x[7:6],x1[7:6]);
recursive_stage1 s03(x[7:6],x[9:8],x1[9:8]);
recursive_stage1 s04(x[9:8],x[11:10],x1[11:10]);
recursive_stage1 s05(x[11:10],x[13:12],x1[13:12]);
recursive_stage1 s06(x[13:12],x[15:14],x1[15:14]);
recursive_stage1 s07(x[15:14],x[17:16],x1[17:16]);
recursive_stage1 s08(x[17:16],x[19:18],x1[19:18]);
recursive_stage1 s09(x[19:18],x[21:20],x1[21:20]);
recursive_stage1 s10(x[21:20],x[23:22],x1[23:22]);
recursive_stage1 s11(x[23:22],x[25:24],x1[25:24]);
recursive_stage1 s12(x[25:24],x[27:26],x1[27:26]);
recursive_stage1 s13(x[27:26],x[29:28],x1[29:28]);
recursive_stage1 s14(x[29:28],x[31:30],x1[31:30]);
recursive_stage1 s15(x[31:30],x[33:32],x1[33:32]);
recursive_stage1 s16(x[33:32],x[35:34],x1[35:34]);
recursive_stage1 s17(x[35:34],x[37:36],x1[37:36]);
recursive_stage1 s18(x[37:36],x[39:38],x1[39:38]);
recursive_stage1 s19(x[39:38],x[41:40],x1[41:40]);
recursive_stage1 s20(x[41:40],x[43:42],x1[43:42]);
recursive_stage1 s21(x[43:42],x[45:44],x1[45:44]);
recursive_stage1 s22(x[45:44],x[47:46],x1[47:46]);
recursive_stage1 s23(x[47:46],x[49:48],x1[49:48]);

wire [49:0] x2;  //recursive doubling stage2
assign x2[3:0]=x1[3:0];

recursive_stage1 s101(x1[1:0],x1[5:4],x2[5:4]);
recursive_stage1 s102(x1[3:2],x1[7:6],x2[7:6]);
recursive_stage1 s103(x1[5:4],x1[9:8],x2[9:8]);
recursive_stage1 s104(x1[7:6],x1[11:10],x2[11:10]);
recursive_stage1 s105(x1[9:8],x1[13:12],x2[13:12]);
recursive_stage1 s106(x1[11:10],x1[15:14],x2[15:14]);
recursive_stage1 s107(x1[13:12],x1[17:16],x2[17:16]);
recursive_stage1 s108(x1[15:14],x1[19:18],x2[19:18]);
recursive_stage1 s109(x1[17:16],x1[21:20],x2[21:20]);
recursive_stage1 s110(x1[19:18],x1[23:22],x2[23:22]);
recursive_stage1 s111(x1[21:20],x1[25:24],x2[25:24]);
recursive_stage1 s112(x1[23:22],x1[27:26],x2[27:26]);
recursive_stage1 s113(x1[25:24],x1[29:28],x2[29:28]);
recursive_stage1 s114(x1[27:26],x1[31:30],x2[31:30]);
recursive_stage1 s115(x1[29:28],x1[33:32],x2[33:32]);
recursive_stage1 s116(x1[31:30],x1[35:34],x2[35:34]);
recursive_stage1 s117(x1[33:32],x1[37:36],x2[37:36]);
recursive_stage1 s118(x1[35:34],x1[39:38],x2[39:38]);
recursive_stage1 s119(x1[37:36],x1[41:40],x2[41:40]);
recursive_stage1 s120(x1[39:38],x1[43:42],x2[43:42]);
recursive_stage1 s121(x1[41:40],x1[45:44],x2[45:44]);
recursive_stage1 s122(x1[43:42],x1[47:46],x2[47:46]);
recursive_stage1 s123(x1[45:44],x1[49:48],x2[49:48]);

wire [49:0] x3;  //recursive doubling stage3
assign x3[7:0]=x2[7:0];

recursive_stage1 s203(x2[1:0],x2[9:8],x3[9:8]);
recursive_stage1 s204(x2[3:2],x2[11:10],x3[11:10]);
recursive_stage1 s205(x2[5:4],x2[13:12],x3[13:12]);
recursive_stage1 s206(x2[7:6],x2[15:14],x3[15:14]);
recursive_stage1 s207(x2[9:8],x2[17:16],x3[17:16]);
recursive_stage1 s208(x2[11:10],x2[19:18],x3[19:18]);
recursive_stage1 s209(x2[13:12],x2[21:20],x3[21:20]);
recursive_stage1 s210(x2[15:14],x2[23:22],x3[23:22]);
recursive_stage1 s211(x2[17:16],x2[25:24],x3[25:24]);
recursive_stage1 s212(x2[19:18],x2[27:26],x3[27:26]);
recursive_stage1 s213(x2[21:20],x2[29:28],x3[29:28]);
recursive_stage1 s214(x2[23:22],x2[31:30],x3[31:30]);
recursive_stage1 s215(x2[25:24],x2[33:32],x3[33:32]);
recursive_stage1 s216(x2[27:26],x2[35:34],x3[35:34]);
recursive_stage1 s217(x2[29:28],x2[37:36],x3[37:36]);
recursive_stage1 s218(x2[31:30],x2[39:38],x3[39:38]);
recursive_stage1 s219(x2[33:32],x2[41:40],x3[41:40]);
recursive_stage1 s220(x2[35:34],x2[43:42],x3[43:42]);
recursive_stage1 s221(x2[37:36],x2[45:44],x3[45:44]);
recursive_stage1 s222(x2[39:38],x2[47:46],x3[47:46]);
recursive_stage1 s223(x2[41:40],x2[49:48],x3[49:48]);

wire [49:0] x4;  //recursive doubling stage 4
assign x4[15:0]=x3[15:0];

recursive_stage1 s307(x3[1:0],x3[17:16],x4[17:16]);
recursive_stage1 s308(x3[3:2],x3[19:18],x4[19:18]);
recursive_stage1 s309(x3[5:4],x3[21:20],x4[21:20]);
recursive_stage1 s310(x3[7:6],x3[23:22],x4[23:22]);
recursive_stage1 s311(x3[9:8],x3[25:24],x4[25:24]);
recursive_stage1 s312(x3[11:10],x3[27:26],x4[27:26]);
recursive_stage1 s313(x3[13:12],x3[29:28],x4[29:28]);
recursive_stage1 s314(x3[15:14],x3[31:30],x4[31:30]);
recursive_stage1 s315(x3[17:16],x3[33:32],x4[33:32]);
recursive_stage1 s316(x3[19:18],x3[35:34],x4[35:34]);
recursive_stage1 s317(x3[21:20],x3[37:36],x4[37:36]);
recursive_stage1 s318(x3[23:22],x3[39:38],x4[39:38]);
recursive_stage1 s319(x3[25:24],x3[41:40],x4[41:40]);
recursive_stage1 s320(x3[27:26],x3[43:42],x4[43:42]);
recursive_stage1 s321(x3[29:28],x3[45:44],x4[45:44]);
recursive_stage1 s322(x3[31:30],x3[47:46],x4[47:46]);
recursive_stage1 s323(x3[33:32],x3[49:48],x4[49:48]);

wire [49:0] x5;  //recursive doubling stage 5
assign x5[31:0]=x4[31:0];

recursive_stage1 s415(x4[1:0],x4[33:32],x5[33:32]);
recursive_stage1 s416(x4[3:2],x4[35:34],x5[35:34]);
recursive_stage1 s417(x4[5:4],x4[37:36],x5[37:36]);
recursive_stage1 s418(x4[7:6],x4[39:38],x5[39:38]);
recursive_stage1 s419(x4[9:8],x4[41:40],x5[41:40]);
recursive_stage1 s420(x4[11:10],x4[43:42],x5[43:42]);
recursive_stage1 s421(x4[13:12],x4[45:44],x5[45:44]);
recursive_stage1 s422(x4[15:14],x4[47:46],x5[47:46]);
recursive_stage1 s423(x4[17:16],x4[49:48],x5[49:48]);

 // final sum and carry

assign sum[0]=a[0]^b[0]^x5[0];
assign sum[1]=a[1]^b[1]^x5[2];
assign sum[2]=a[2]^b[2]^x5[4];
assign sum[3]=a[3]^b[3]^x5[6];
assign sum[4]=a[4]^b[4]^x5[8];
assign sum[5]=a[5]^b[5]^x5[10];
assign sum[6]=a[6]^b[6]^x5[12];
assign sum[7]=a[7]^b[7]^x5[14];
assign sum[8]=a[8]^b[8]^x5[16];
assign sum[9]=a[9]^b[9]^x5[18];
assign sum[10]=a[10]^b[10]^x5[20];
assign sum[11]=a[11]^b[11]^x5[22];
assign sum[12]=a[12]^b[12]^x5[24];
assign sum[13]=a[13]^b[13]^x5[26];
assign sum[14]=a[14]^b[14]^x5[28];
assign sum[15]=a[15]^b[15]^x5[30];
assign sum[16]=a[16]^b[16]^x5[32];
assign sum[17]=a[17]^b[17]^x5[34];
assign sum[18]=a[18]^b[18]^x5[36];
assign sum[19]=a[19]^b[19]^x5[38];
assign sum[20]=a[20]^b[20]^x5[40];
assign sum[21]=a[21]^b[21]^x5[42];
assign sum[22]=a[22]^b[22]^x5[44];
assign sum[23]=a[23]^b[23]^x5[46];

kgp_carry kkc(x[49:48],x5[47:46],carry);

endmodule



//mux31to1

module mux32to1_24(out,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,s4,s3,s2,s1,s0);
input [23:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31;
input s4,s3,s2,s1,s0;
output [23:0] out;

//level 1 

reg [23:0] out;

always@(i0 or i1 or i2 or i3 or i4 or i5 or i6 or i7 or i8 or i9 or i10 or i11 or i12 or i13 or i14 or i15 or i16 or i17 or i18 or i19 or i20 or i21 or i22 or i23 or i24 or i25 or i26 or i27 or i28 or i29 or i30 or i31 or s4 or s3 or s2 or s1 or s0)
begin 
case({s4,s3,s2,s1,s0})
5'b00000: out = i0;
5'b00001: out = i1;
5'b00010: out = i2;
5'b00011: out = i3;
5'b00100: out = i4;
5'b00101: out = i5;
5'b00110: out = i6;
5'b00111: out = i7;
5'b01000: out = i8;
5'b01001: out = i9;
5'b01010: out = i10;
5'b01011: out = i11;
5'b01100: out = i12;
5'b01101: out = i13;
5'b01110: out = i14;
5'b01111: out = i15;
5'b10000: out = i16;
5'b10001: out = i17;
5'b10010: out = i18;
5'b10011: out = i19;
5'b10100: out = i20;
5'b10101: out = i21;
5'b10110: out = i22;
5'b10111: out = i23;
5'b11000: out = i24;
5'b11001: out = i25;
5'b11010: out = i26;
5'b11011: out = i27;
5'b11100: out = i28;
5'b11101: out = i29;
5'b11110: out = i30;
5'b11111: out = i31;
default: out = 1'bx;
endcase
end 


endmodule


//mux16to1

module mux16to1_24(o,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,s);

input [23:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15;
input [3:0] s;
output [23:0] o;
reg [23:0] o;

always@(i0 or i1 or i2 or i3 or i4 or i5 or i6 or i7 or i8 or i9 or i10 or i11 or i12 or i13 or i14 or i15 or s)
	begin
		case(s)
		 4'b0000:o=i0;
		 4'b0001:o=i1;
		 4'b0010:o=i2;
		 4'b0011:o=i3;
		 4'b0100:o=i4;
		 4'b0101:o=i5;
		 4'b0110:o=i6;
		 4'b0111:o=i7;
		 4'b1000:o=i8;
		 4'b1001:o=i9;
		 4'b1010:o=i10;
		 4'b1011:o=i11;
		 4'b1100:o=i12;
		 4'b1101:o=i13;
		 4'b1110:o=i14;
		 4'b1111:o=i15;
		 //default:o=1'bx;
		endcase
	end



endmodule




//mux8to1

module mux8to1_24(o,i0,i1,i2,i3,i4,i5,i6,i7,s);

input [23:0] i0,i1,i2,i3,i4,i5,i6,i7;
input [2:0] s;
output [23:0] o;
reg [23:0] o;

always@(i0 or i1 or i2 or i3 or i4 or i5 or i6 or i7 or s)
	begin
		case(s)
		 3'b000:o=i0;
		 3'b001:o=i1;
		 3'b010:o=i2;
		 3'b011:o=i3;
		 3'b100:o=i4;
		 3'b101:o=i5;
		 3'b110:o=i6;
		 3'b111:o=i7;
		 //default:o=1'bx;
		endcase
	end


endmodule


//mux4to1

module mux4to1_24(y,in0,in1,in2,in3,sel);

input [23:0] in0,in1,in2,in3;
input [1:0] sel;
output [23:0] y;

reg [23:0] y;
always@(in0 or in1 or in2 or in3 or sel)
begin
case(sel)
2'b00:y=in0;  
2'b01:y=in1;
2'b10:y=in2;	
2'b11:y=in3;  
//default:y=1'bx;
endcase   
end


endmodule



//2 to 1 multiplexer design

module mux2to1_24(out,i1,i2,s);

input [23:0] i1,i2;
input s;
output [23:0] out;
reg [23:0] out;

always@(i1 or i2 or s)
	begin
	 case(s)
	  1'b0:out=i1;
	  1'b1:out=i2;
	 endcase
	end

endmodule


//mux5 to 1

module mux5to1_24(o,o1,o2,o3,o4,o5,dir);

input [2:0] dir;
input [23:0] o1,o2,o3,o4,o5;
output [23:0] o;

reg [23:0] o;

always@(o1 or o2 or o3 or o4 or o5 or dir)
	begin
	 case(dir)
	  3'b000: o=o1;
	  3'b001: o=o2;
	  3'b010: o=o3;
	  3'b011: o=o4;
	  3'b100: o=o5;	  
	default: o = 1'bx;
	 endcase
	end

endmodule


//mux32to1

module mux32to1_1(out,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,s4,s3,s2,s1,s0);
input i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31,s4,s3,s2,s1,s0;
output out;

//level 1 

reg out;

always@(i0 or i1 or i2 or i3 or i4 or i5 or i6 or i7 or i8 or i9 or i10 or i11 or i12 or i13 or i14 or i15 or i16 or i17 or i18 or i19 or i20 or i21 or i22 or i23 or i24 or i25 or i26 or i27 or i28 or i29 or i30 or i31 or s4 or s3 or s2 or s1 or s0)
begin 
case({s4,s3,s2,s1,s0})
5'b00000: out = i0;
5'b00001: out = i1;
5'b00010: out = i2;
5'b00011: out = i3;
5'b00100: out = i4;
5'b00101: out = i5;
5'b00110: out = i6;
5'b00111: out = i7;
5'b01000: out = i8;
5'b01001: out = i9;
5'b01010: out = i10;
5'b01011: out = i11;
5'b01100: out = i12;
5'b01101: out = i13;
5'b01110: out = i14;
5'b01111: out = i15;
5'b10000: out = i16;
5'b10001: out = i17;
5'b10010: out = i18;
5'b10011: out = i19;
5'b10100: out = i20;
5'b10101: out = i21;
5'b10110: out = i22;
5'b10111: out = i23;
5'b11000: out = i24;
5'b11001: out = i25;
5'b11010: out = i26;
5'b11011: out = i27;
5'b11100: out = i28;
5'b11101: out = i29;
5'b11110: out = i30;
5'b11111: out = i31;
default: out = 1'bx;
endcase
end 


endmodule


//mux16to1

module mux16to1_1(o,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,s);

input i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15;
input [3:0] s;
output o;
reg o;

always@(i0 or i1 or i2 or i3 or i4 or i5 or i6 or i7 or i8 or i9 or i10 or i11 or i12 or i13 or i14 or i15 or s)
	begin
		case(s)
		 4'b0000:o=i0;
		 4'b0001:o=i1;
		 4'b0010:o=i2;
		 4'b0011:o=i3;
		 4'b0100:o=i4;
		 4'b0101:o=i5;
		 4'b0110:o=i6;
		 4'b0111:o=i7;
		 4'b1000:o=i8;
		 4'b1001:o=i9;
		 4'b1010:o=i10;
		 4'b1011:o=i11;
		 4'b1100:o=i12;
		 4'b1101:o=i13;
		 4'b1110:o=i14;
		 4'b1111:o=i15;
		 //default:o=1'bx;
		endcase
	end


endmodule


//mux8to1

module mux8to1_1(o,i0,i1,i2,i3,i4,i5,i6,i7,s);

input i0,i1,i2,i3,i4,i5,i6,i7;
input [2:0] s;
output o;
reg o;

always@(i0 or i1 or i2 or i3 or i4 or i5 or i6 or i7 or s)
	begin
		case(s)
		 3'b000:o=i0;
		 3'b001:o=i1;
		 3'b010:o=i2;
		 3'b011:o=i3;
		 3'b100:o=i4;
		 3'b101:o=i5;
		 3'b110:o=i6;
		 3'b111:o=i7;
		 //default:o=1'bx;
		endcase
	end


endmodule


//mux4to1

module mux4to1_1(y,in0,in1,in2,in3,sel);

input in0,in1,in2,in3;
input [1:0] sel;
output y;

reg y;
always@(in0 or in1 or in2 or in3 or sel)
begin
case(sel)
2'b00:y=in0;  
2'b01:y=in1;
2'b10:y=in2;	
2'b11:y=in3;  
//default:y=1'bx;
endcase   
end

endmodule


//2 to 1 multiplexer design

module mux2to1_1(out,i1,i2,s);

input i1,i2,s;
output out;
reg out;

always@(i1 or i2 or s)
	begin
	 case(s)
	  1'b0:out=i1;
	  1'b1:out=i2;
	 endcase
	end

endmodule


//mux5 to 1

module mux5to1_1(o,o1,o2,o3,o4,o5,dir);

input [2:0] dir;
input o1,o2,o3,o4,o5;
output o;

reg o;

always@(o1 or o2 or o3 or o4 or o5 or dir)
	begin
	 case(dir)
	  3'b000: o=o1;
	  3'b001: o=o2;
	  3'b010: o=o3;
	  3'b011: o=o4;
	  3'b100: o=o5;
	  
	default: o = 1'bx;
	 endcase
	end

endmodule



















































`default_nettype wire
